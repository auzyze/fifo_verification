class Environment;

  Generator     gen;
  
  mailbox       gen2drv;
  mailbox       drv2scb;
  mailbox       mon2scb;
  
  event         drv2gen;
  
  Driver        drv;
  Monitor       mon;
  Scoreboard    scb;
  Coverage      cov;
  
  Config        cfg;          //used to configure TB
  
  CPU_driver    cpu;          //driver used to configure DUT

  vFifo_TB      test_intf;    //virtual interface
  vCPU_T        cfg_intf;     //virtual interface
  
  extern function new(input vFifo_TB  test_intf,
                      input vCPU_T    cfg_intf
                      );
  
  extern virtual function void gen_cfg();
  extern virtual function void build();
  extern virtual task run();
  extern virtual function void wrap_up();
  
endclass: Environment

///////////////////////////////////////////////////
//construct an environment instance
function Environment::new(input vFifo_TB  test_intf,
                          input vCPU_T    cfg_intf
                          );
  this.test_intf = test_intf;
  this.cfg_intf = cfg_intf;  
  cfg = new();
endfunction : new
  

///////////////////////////////////////////////////
//configure ??
function void Environment::gen_cfg();
  assert(cfg.randomize());
  cfg.display();
endfunction : gen_cfg


//////////////////////////////////////////////////
//Build the environment objects
function void Environment::build();
  cpu = new(cfg_intf,cfg);            //construct CPU driver with cfg info
  gen = new();
  drv = new();
  
  gen2drv = new();                    //mailbox X 3
  drv2scb = new();
  mon2scb = new();
  
  drv2gen = new();                    //event
  
  scb = new(cfg);                     //construct scoreboard with cfg info
  cov = new();
  mon = new();  
  
endfunction : build


//////////////////////////////////////////////////////
//Start the transactors: generator, driver, monior
task Environment::run();
  
  //The CPU interface initializes before anyone else
  cpu.run();
  
  //Generator and Driver
  gen.run();
  drv.run();
  
  //Monitor
  mon.run();
  
  //wait for data to flow through DUT, monitor and scoreboard
  repeat (10000)@(test_intf.cb);
  
endtask : run
  
  
  
///////////////////////////////////////////
//Post-run cleanup / reporting
function void Environment::wrap_up();
  $display("@%0t: End of sim, %0d errors, %0d warnings",
            $time, cfg.nErrors, cfg.nWarnings);
  scb.wrap_up;
endfunction : wrap_up



////////////////////////////////////////////////
//Define basic transaction : single write or read
class fifo_op;
  rand bit [1:0]  op_type;
  rand bit [15:0] op_len;
  
  rand bit [31:0] data [];
    
  bit [31:0] rd_data;
  bit full;
  bit empty;
  bit afull;
  bit aempty;

  //static bit [15:0] wr_count;
  //static bit [15:0] rd_count;

  //extern function new();
  //extern function void post_randomize();
    
endclass : fifo_op



///////////////////////////////////////////////////////
///////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////
//FIFO Operation Generator
class Generator;
  fifo_op gen_op;
  mailbox gen2drv;
  event   drv2gen;
  
  int     op_num;
  
  function new(input mailbox gen2drv,
               input event drv2gen,
               input int op_num);
    this.gen2drv = gen2drv;
    this.drv2gen = drv2gen;
    this.op_num = op_num;
    gen_op = new();
  endfunction : new
  
  task run();
    repeat (op_num) begin
      assert (gen_op.randomize());
      gen2drv.put(gen_op);
      @drv2gen; //Wait for driver to finish with it
    end
  endtask : run
  
endclass : Generator



//////////////////////////////////////////////////////
////////////////////////////////////////////////////////
//Driver
class Driver;
  mailbox gen2drv;
  mailbox drv2scb;
  event   drv2gen;
  vFifo_TB test_intf;     //virtual interface for operation transimitting
  
  extern function new(input mailbox gen2drv,
                      input mailbox drv2scb,
                      input event drv2gen,
                      input vFifo_TB test_intf);
  extern task run();
  extern task send (input fifo_op gen_op);
  
endclass : Driver

//
function Driver::new(input mailbox gen2drv,
                     input event drv2gen,
                     input vFifo_TB test_intf);
  this.gen2drv = gen2drv;
  this.drv2gen = drv2gen;
  this.test_intf = test_intf;
endfunction : new

//run() : run the driver
task Driver::run();
  fifo_op gen_op;
  
  //Initialize ports
  test_intf.cb.wr_en <= 0;
  test_intf.cb.wr_data <= 0;
  test_intf.cb.rd_en <= 0;
  
  forever begin
    gen2drv.peek(gen_op);      //"peek" task gets a copy of data in mailbox but doesn't remove it
    send(gen_op);
    gen2drv.get(gen_op);       //remove the data with "get" task after operation has been sent
    ->drv2gen;
  end
endtask : run

//send() : Send a operation into DUT
task Driver::send(input fifo_op gen_op);
  for (i=0; i<gen_op.op_len; i++) begin
    case (op_type)
      2'b00:
        test_intf.wr_en <= 0;
        test_intf.rd_en <= 0;
        test_intf.wr_data <= 0;
      2'b01:
        test_intf.wr_en <= 0;
        test_intf.rd_en <= 1;
        test_intf.wr_data <= 0;      
      2'b10:
        test_intf.wr_en <= 1;
        test_intf.rd_en <= 0;
        test_intf.wr_data <= gen_op.wr_data[];  // ?????        
      2'b11:
        test_intf.wr_en <= 1;
        test_intf.rd_en <= 1;
        test_intf.wr_data <= gen_op.wr_data[];  // ?????        
    endcase
    @test_intf.cb;
  end
  
endtask : Driver



/////////////////////////////////////////////////////////////
//Monitor

class Monitor;
  vFifo_TB op_intf;
  
  extern function new(input vFifo_TB op_intf);
  extern task run();
  extern task receive(output RData output_d);    //what should be received?
endclass : Monitor

//new
function Monitor::new(input vFifo_TB op_intf);
  this.op_intf = op_intf;
endfunction


task Monitor::run();
  RData output_d;
  
  forever begin
    receive(output_d);
  end
  
endtask : run


//receive task
task Monitor::receive(output RData output_d)

.....

endtask : receive



///////////////////////////////////////////////////
//the scoreboard class









